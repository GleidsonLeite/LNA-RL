.title LNA Test
.include /edatools/opentools/skywater-pdk/libraries/sky130_fd_pr/latest/models/corners/tt.spice
.subckt LNA IN OUT VCC VDD VPOL1 VPOL2 GND
.subckt NFET1 DRAIN GATE SOURCE SUBSTRATE
XM1 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 L=2.2 W=68.3 ad='W*0.29' as_='W*0.29' mult=1 nf=1 nrd='0.29/W' nrs='0.29/W' pd='2*(W+0.29)' ps='2*(W+0.29)' sa=0 sb=0 sd=0
.ends NFET1

.subckt PFET2 DRAIN GATE SOURCE SUBSTRATE
XM1 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__pfet_01v8 L=39.9 W=1.1 ad='W*0.29' as_='W*0.29' mult=1 nf=1 nrd='0.29/W' nrs='0.29/W' pd='2*(W+0.29)' ps='2*(W+0.29)' sa=0 sb=0 sd=0
.ends PFET2

.subckt NFET3 DRAIN GATE SOURCE SUBSTRATE
XM1 DRAIN GATE SOURCE SUBSTRATE sky130_fd_pr__nfet_01v8 L=48 W=6.5 ad='W*0.29' as_='W*0.29' mult=1 nf=1 nrd='0.29/W' nrs='0.29/W' pd='2*(W+0.29)' ps='2*(W+0.29)' sa=0 sb=0 sd=0
.ends NFET3
LLG IN PLG 5.8e-09
RRPOL1 PLG VPOL1 19939
XM1 PRF PLG GND GND NFETW1
CC1 PC1 PLG 1.97e-11
RRF PC1 PRF 19540
XM2 VCC PC1 PRF GND PFET2
CCDEC VCC GND 1e-06
CCM1 PRF PCM1 4.7e-12
RRPOL2 PCM1 VPOL2 13548
XM3 PM3 PCM1 GND GND NFETW3
LLPK VDD PM3 7.6e-09
CCM2 PM3 OUT 6.5e-13
CCM3 PM3 GND 4.7e-12
.ends LNA

.subckt SourceCircuit IN VCC VDD VPOL1 VPOL2 GND
Vsignal IN GND DC 0.5V AC 1V SIN(0V 1V 50Hz 0s 0Hz)
VVCC VCC GND 1.8
VVDD VDD GND 1.8
VVPOL1 VPOL1 GND 1.1
VVPOL2 VPOL2 GND 0.68
.ends SourceCircuit
Xamplifier IN OUT VCC VDD VPOL1 VPOL2 0 LNA
Xsource IN VCC VDD VPOL1 VPOL2 0 SourceCircuit
RRtest OUT 0 50